`timescale 1ns / 1ps

module rom_sign_mag_adder(
    input wire clk,
    input wire [3:0] a, b,
    output wire [3:0] data
    );
    
    reg [3:0] rom_data, data_reg;
    
    always @(posedge clk)
        data_reg <= rom_data;
        
    always @*
        case({a,b})
            8'b11111111: rom_data=4'b0000;
            8'b11111110: rom_data=4'b0000;
            8'b11111101: rom_data=4'b0000;
            8'b11111100: rom_data=4'b0000;
            8'b11111011: rom_data=4'b0000;
            8'b11111010: rom_data=4'b0000;
            8'b11111001: rom_data=4'b0000;
            8'b11110000: rom_data=4'b1111;
            8'b11110001: rom_data=4'b1110;
            8'b11110010: rom_data=4'b1101;
            8'b11110011: rom_data=4'b1100;
            8'b11110100: rom_data=4'b1011;
            8'b11110101: rom_data=4'b1010;
            8'b11110110: rom_data=4'b1001;
            8'b11110111: rom_data=4'b0000;
            8'b11101111: rom_data=4'b0000;
            8'b11101110: rom_data=4'b0000;
            8'b11101101: rom_data=4'b0000;
            8'b11101100: rom_data=4'b0000;
            8'b11101011: rom_data=4'b0000;
            8'b11101010: rom_data=4'b0000;
            8'b11101001: rom_data=4'b1111;
            8'b11100000: rom_data=4'b1110;
            8'b11100001: rom_data=4'b1101;
            8'b11100010: rom_data=4'b1100;
            8'b11100011: rom_data=4'b1011;
            8'b11100100: rom_data=4'b1010;
            8'b11100101: rom_data=4'b1001;
            8'b11100110: rom_data=4'b0000;
            8'b11100111: rom_data=4'b0001;
            8'b11011111: rom_data=4'b0000;
            8'b11011110: rom_data=4'b0000;
            8'b11011101: rom_data=4'b0000;
            8'b11011100: rom_data=4'b0000;
            8'b11011011: rom_data=4'b0000;
            8'b11011010: rom_data=4'b1111;
            8'b11011001: rom_data=4'b1110;
            8'b11010000: rom_data=4'b1101;
            8'b11010001: rom_data=4'b1100;
            8'b11010010: rom_data=4'b1011;
            8'b11010011: rom_data=4'b1010;
            8'b11010100: rom_data=4'b1001;
            8'b11010101: rom_data=4'b0000;
            8'b11010110: rom_data=4'b0001;
            8'b11010111: rom_data=4'b0010;
            8'b11001111: rom_data=4'b0000;
            8'b11001110: rom_data=4'b0000;
            8'b11001101: rom_data=4'b0000;
            8'b11001100: rom_data=4'b0000;
            8'b11001011: rom_data=4'b1111;
            8'b11001010: rom_data=4'b1110;
            8'b11001001: rom_data=4'b1101;
            8'b11000000: rom_data=4'b1100;
            8'b11000001: rom_data=4'b1011;
            8'b11000010: rom_data=4'b1010;
            8'b11000011: rom_data=4'b1001;
            8'b11000100: rom_data=4'b0000;
            8'b11000101: rom_data=4'b0001;
            8'b11000110: rom_data=4'b0010;
            8'b11000111: rom_data=4'b0011;
            8'b10111111: rom_data=4'b0000;
            8'b10111110: rom_data=4'b0000;
            8'b10111101: rom_data=4'b0000;
            8'b10111100: rom_data=4'b1111;
            8'b10111011: rom_data=4'b1110;
            8'b10111010: rom_data=4'b1101;
            8'b10111001: rom_data=4'b1100;
            8'b10110000: rom_data=4'b1011;
            8'b10110001: rom_data=4'b1010;
            8'b10110010: rom_data=4'b1001;
            8'b10110011: rom_data=4'b0000;
            8'b10110100: rom_data=4'b0001;
            8'b10110101: rom_data=4'b0010;
            8'b10110110: rom_data=4'b0011;
            8'b10110111: rom_data=4'b0100;
            8'b10101111: rom_data=4'b0000;
            8'b10101110: rom_data=4'b0000;
            8'b10101101: rom_data=4'b1111;
            8'b10101100: rom_data=4'b1110;
            8'b10101011: rom_data=4'b1101;
            8'b10101010: rom_data=4'b1100;
            8'b10101001: rom_data=4'b1011;
            8'b10100000: rom_data=4'b1010;
            8'b10100001: rom_data=4'b1001;
            8'b10100010: rom_data=4'b0000;
            8'b10100011: rom_data=4'b0001;
            8'b10100100: rom_data=4'b0010;
            8'b10100101: rom_data=4'b0011;
            8'b10100110: rom_data=4'b0100;
            8'b10100111: rom_data=4'b0101;
            8'b10011111: rom_data=4'b0000;
            8'b10011110: rom_data=4'b1111;
            8'b10011101: rom_data=4'b1110;
            8'b10011100: rom_data=4'b1101;
            8'b10011011: rom_data=4'b1100;
            8'b10011010: rom_data=4'b1011;
            8'b10011001: rom_data=4'b1010;
            8'b10010000: rom_data=4'b1001;
            8'b10010001: rom_data=4'b0000;
            8'b10010010: rom_data=4'b0001;
            8'b10010011: rom_data=4'b0010;
            8'b10010100: rom_data=4'b0011;
            8'b10010101: rom_data=4'b0100;
            8'b10010110: rom_data=4'b0101;
            8'b10010111: rom_data=4'b0110;
            8'b00001111: rom_data=4'b1111;
            8'b00001110: rom_data=4'b1110;
            8'b00001101: rom_data=4'b1101;
            8'b00001100: rom_data=4'b1100;
            8'b00001011: rom_data=4'b1011;
            8'b00001010: rom_data=4'b1010;
            8'b00001001: rom_data=4'b1001;
            8'b00000000: rom_data=4'b0000;
            8'b00000001: rom_data=4'b0001;
            8'b00000010: rom_data=4'b0010;
            8'b00000011: rom_data=4'b0011;
            8'b00000100: rom_data=4'b0100;
            8'b00000101: rom_data=4'b0101;
            8'b00000110: rom_data=4'b0110;
            8'b00000111: rom_data=4'b0111;
            8'b00011111: rom_data=4'b1110;
            8'b00011110: rom_data=4'b1101;
            8'b00011101: rom_data=4'b1100;
            8'b00011100: rom_data=4'b1011;
            8'b00011011: rom_data=4'b1010;
            8'b00011010: rom_data=4'b1001;
            8'b00011001: rom_data=4'b0000;
            8'b00010000: rom_data=4'b0001;
            8'b00010001: rom_data=4'b0010;
            8'b00010010: rom_data=4'b0011;
            8'b00010011: rom_data=4'b0100;
            8'b00010100: rom_data=4'b0101;
            8'b00010101: rom_data=4'b0110;
            8'b00010110: rom_data=4'b0111;
            8'b00010111: rom_data=4'b0000;
            8'b00101111: rom_data=4'b1101;
            8'b00101110: rom_data=4'b1100;
            8'b00101101: rom_data=4'b1011;
            8'b00101100: rom_data=4'b1010;
            8'b00101011: rom_data=4'b1001;
            8'b00101010: rom_data=4'b0000;
            8'b00101001: rom_data=4'b0001;
            8'b00100000: rom_data=4'b0010;
            8'b00100001: rom_data=4'b0011;
            8'b00100010: rom_data=4'b0100;
            8'b00100011: rom_data=4'b0101;
            8'b00100100: rom_data=4'b0110;
            8'b00100101: rom_data=4'b0111;
            8'b00100110: rom_data=4'b0000;
            8'b00100111: rom_data=4'b0000;
            8'b00111111: rom_data=4'b1100;
            8'b00111110: rom_data=4'b1011;
            8'b00111101: rom_data=4'b1010;
            8'b00111100: rom_data=4'b1001;
            8'b00111011: rom_data=4'b0000;
            8'b00111010: rom_data=4'b0001;
            8'b00111001: rom_data=4'b0010;
            8'b00110000: rom_data=4'b0011;
            8'b00110001: rom_data=4'b0100;
            8'b00110010: rom_data=4'b0101;
            8'b00110011: rom_data=4'b0110;
            8'b00110100: rom_data=4'b0111;
            8'b00110101: rom_data=4'b0000;
            8'b00110110: rom_data=4'b0000;
            8'b00110111: rom_data=4'b0000;
            8'b01001111: rom_data=4'b1011;
            8'b01001110: rom_data=4'b1010;
            8'b01001101: rom_data=4'b1001;
            8'b01001100: rom_data=4'b0000;
            8'b01001011: rom_data=4'b0001;
            8'b01001010: rom_data=4'b0010;
            8'b01001001: rom_data=4'b0011;
            8'b01000000: rom_data=4'b0100;
            8'b01000001: rom_data=4'b0101;
            8'b01000010: rom_data=4'b0110;
            8'b01000011: rom_data=4'b0111;
            8'b01000100: rom_data=4'b0000;
            8'b01000101: rom_data=4'b0000;
            8'b01000110: rom_data=4'b0000;
            8'b01000111: rom_data=4'b0000;
            8'b01011111: rom_data=4'b1010;
            8'b01011110: rom_data=4'b1001;
            8'b01011101: rom_data=4'b0000;
            8'b01011100: rom_data=4'b0001;
            8'b01011011: rom_data=4'b0010;
            8'b01011010: rom_data=4'b0011;
            8'b01011001: rom_data=4'b0100;
            8'b01010000: rom_data=4'b0101;
            8'b01010001: rom_data=4'b0110;
            8'b01010010: rom_data=4'b0111;
            8'b01010011: rom_data=4'b0000;
            8'b01010100: rom_data=4'b0000;
            8'b01010101: rom_data=4'b0000;
            8'b01010110: rom_data=4'b0000;
            8'b01010111: rom_data=4'b0000;
            8'b01101111: rom_data=4'b1001;
            8'b01101110: rom_data=4'b0000;
            8'b01101101: rom_data=4'b0001;
            8'b01101100: rom_data=4'b0010;
            8'b01101011: rom_data=4'b0011;
            8'b01101010: rom_data=4'b0100;
            8'b01101001: rom_data=4'b0101;
            8'b01100000: rom_data=4'b0110;
            8'b01100001: rom_data=4'b0111;
            8'b01100010: rom_data=4'b0000;
            8'b01100011: rom_data=4'b0000;
            8'b01100100: rom_data=4'b0000;
            8'b01100101: rom_data=4'b0000;
            8'b01100110: rom_data=4'b0000;
            8'b01100111: rom_data=4'b0000;
            8'b01111111: rom_data=4'b0000;
            8'b01111110: rom_data=4'b0001;
            8'b01111101: rom_data=4'b0010;
            8'b01111100: rom_data=4'b0011;
            8'b01111011: rom_data=4'b0100;
            8'b01111010: rom_data=4'b0101;
            8'b01111001: rom_data=4'b0110;
            8'b01110000: rom_data=4'b0111;
            8'b01110001: rom_data=4'b0000;
            8'b01110010: rom_data=4'b0000;
            8'b01110011: rom_data=4'b0000;
            8'b01110100: rom_data=4'b0000;
            8'b01110101: rom_data=4'b0000;
            8'b01110110: rom_data=4'b0000;
            8'b01110111: rom_data=4'b0000;
        endcase
   
    assign data = data_reg; 
endmodule
